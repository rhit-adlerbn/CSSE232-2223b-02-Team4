module tb_InstMem

endmodule 