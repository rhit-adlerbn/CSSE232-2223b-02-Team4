module REG

endmodule 