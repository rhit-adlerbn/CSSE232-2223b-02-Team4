module tb_ImmGen

endmodule 