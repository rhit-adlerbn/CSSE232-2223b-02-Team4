module IMMGEN

endmodule 