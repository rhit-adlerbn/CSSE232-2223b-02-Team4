module ALU

endmodule 