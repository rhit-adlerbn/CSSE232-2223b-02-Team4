module tb_Reg

endmodule 