module tb_Alu

endmodule 