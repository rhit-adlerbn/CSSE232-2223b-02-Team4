module tb_DataMem

endmodule 