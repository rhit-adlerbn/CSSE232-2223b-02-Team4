module PC

endmodule