module DoomProcessor

endmodule
