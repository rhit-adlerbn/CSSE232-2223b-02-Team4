module tb_Pc

endmodule 