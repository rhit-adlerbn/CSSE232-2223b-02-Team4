module INSTMEM

endmodule 