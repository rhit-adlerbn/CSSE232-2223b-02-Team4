module DATAMEM

endmodule 